
package axi_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "axi_seq_item.sv"
    `include "axi_driver.sv"
    `include "axi_monitor.sv"
    `include "axi_agent.sv"
    `include "axi_scoreboard.sv"
    `include "axi_base_seq.sv"

endpackage
